//------------------------------------------------------------
//   Copyright 2010-2019 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------

package spi_virtual_seq_lib_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

import apb_agent_pkg::*;
import spi_agent_pkg::*;
import spi_env_pkg::*;
import spi_bus_sequence_lib_pkg::*;
import spi_sequence_lib_pkg::*;

typedef class spi_vseq_base;
typedef class config_interrupt_vseq;
typedef class config_polling_vseq;
typedef class reg_test_vseq;

`include "top_virtual_seqs/spi_vseq_base.svh"
`include "top_virtual_seqs/config_interrupt_vseq.svh"
`include "top_virtual_seqs/config_polling_vseq.svh"
`include "top_virtual_seqs/reg_test_vseq.svh"



endpackage:spi_virtual_seq_lib_pkg
