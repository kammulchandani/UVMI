/***********************************************************************
 * Testbench top for "dual-top" example for UVM Intermediate lab 1 DMA
 ***********************************************************************
 * Copyright 2019 Mentor Graphics Corporation
 * All Rights Reserved Worldwide
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *       http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or
 * implied.  See the License for the specific language governing
 * permissions and limitations under the License.
 **********************************************************************/

module top_hdl();
  import uvm_pkg::*;

  dma_ifc  dma_if();
  dma_ctrl dma0(dma_if);
  initial begin
    $timeformat(-9,0,"ns",6);
    uvm_config_db #(virtual dma_ifc)::set(null, "uvm_test_top", "dma_if", dma_if);
  end
endmodule
